
module HELLOWORLD (
	clk_clk);	

	input		clk_clk;
endmodule


module HELLO (
	clk_clk);	

	input		clk_clk;
endmodule
